LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ULA1BIT IS
	PORT(x: IN BIT;
		z: OUT BIT);
END ULA1BIT;

ARCHITECTURE logica1 OF ULA1BIT IS
	BEGIN
END logica1;
