LIBRARY ieee, components;
USE ieee.std_logic_1164.all, components.all;

ENTITY ULA1BIT IS
	PORT(x,y: IN BIT;
		z: OUT BIT);
END ULA1BIT;

ARCHITECTURE logica1 OF ULA1BIT IS
	BEGIN
END logica1;
