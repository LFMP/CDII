LIBRARY components;
USE components.all;

ENTITY ULA1BIT IS
	PORT(x,y: IN BIT;
		z: OUT BIT);
END ULA1BIT;

ARCHITECTURE logica1 OF ULA1BIT IS
	BEGIN
END logica1;
